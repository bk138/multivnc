"NSLocalNetworkUsageDescription" = "MultiVNC kräver åtkomst till ditt lokala nätverk för att kunna upptäcka och ansluta till VNC-servrar för fjärrstyrning av skrivbordet.";
